package alu_pkg;
	  import std::*; // some package issue 
	`include "transaction.sv"
	`include "generator.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "reference.sv"	
	`include "scoreboard.sv"
	`include "environment.sv"
	`include "test.sv"
endpackage
