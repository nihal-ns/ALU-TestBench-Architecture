`include "defines.sv"

class monitor;
	transaction trans;
	mailbox #(transaction) mon2scb;
	virtual intf.MONITOR vif;

	function new(mailbox #(transaction) mon2scb, virtual intf.MONITOR vif);
		this.mon2scb = mon2scb;
		this.vif = vif;
	endfunction

	task start();
		repeat(2) @(vif.mon_cb);  // changed to 1
		for(int i=0; i<`no_trans; i++) begin
			trans = new;
			repeat(3) @(vif.mon_cb) // changed 2
			if(vif.mon_cb.MODE && vif.mon_cb.CMD ==9) 
				repeat(1)@(vif.mon_cb);
				
			        /* if(((vif.mon_cb.MODE) && (vif.mon_cb.CMD < 4 || vif.mon_cb.CMD > 7) && (vif.mon_cb.CMD <11)) || ((!vif.mon_cb.MODE) && (vif.mon_cb.CMD < 6 || vif.mon_cb.CMD > 11 ) && (vif.mon_cb.CMD < 14)) && vif.mon_cb.INP_VALID != 2'b11) begin */  
					/* for(int i =0;i<16;i++) begin */ 
						/* @(vif.mon_cb); */
						/* if(i==15) begin */
							/* if(vif.mon_cb.INP_VALID == 2'b11) */
								/* break; */
						/* else */
							/* if(vif.mon_cb.INP_VALID == 2'b11); */
							/* break; */
						/* end */
					/* end */
				/* end */


			/* begin */
				trans.RES = vif.mon_cb.RES;
				trans.OFLOW = vif.mon_cb.OFLOW;
				trans.COUT = vif.mon_cb.COUT;
				trans.E = vif.mon_cb.E;
				trans.G = vif.mon_cb.G;
				trans.L = vif.mon_cb.L;
				trans.ERR = vif.mon_cb.ERR;
				trans.MODE = vif.mon_cb.MODE;
				trans.CMD = vif.mon_cb.CMD;
				trans.OPA = vif.mon_cb.OPA;
				trans.OPB = vif.mon_cb.OPB;
			/* end */
			/* $display("-------------------------------------|| MONITOR ||----------------------------------------------"); */
			if(trans.MODE)
				$display("\n%0t || MONITOR Arithmetic: \t|||cmd:%0d |A:%0d |B:%0d |valid:%0b \n\t\t\t\t|||result:%0d |overflow:%0b |cout:%0b |EGL:%0b%0b%0b |error:%b",$time,trans.CMD,trans.OPA,trans.OPB, trans.INP_VALID, trans.RES, trans.OFLOW, trans.COUT, trans.E, trans.G, trans.L, trans.ERR);
			else
				$display("\n%0t || MONITOR Logical:	|||cmd:%0d |A:%0b |B:%0b |valid:%0b \n\t\t\t\t|||result:%0b |overflow:%0b |cout:%0b |EGL:%0b%0b%0b |error:%0b",$time,trans.CMD,trans.OPA,trans.OPB, trans.INP_VALID, trans.RES, trans.OFLOW, trans.COUT, trans.E, trans.G, trans.L, trans.ERR);
			mon2scb.put(trans);
			//repeat(2)@(vif.mon_cb); 
		end
	endtask
endclass


